library IEEE;
use IEEE.std_logic_1164.all;
--------------------------------------------------------------------------------
package lfsr is

    ----------------------------------------------------------------------------
    -- Types & Constants
    ----------------------------------------------------------------------------
    constant C_TAPTABLE_WIDTH : natural := 5;
    constant C_TAPTABLE_MIN   : natural := 3;
    constant C_TAPTABLE_MAX   : natural := 168;
    type t_taptable is array(C_TAPTABLE_MIN to C_TAPTABLE_MAX, 0 to C_TAPTABLE_WIDTH-1) of natural;

    -- Xilinx XAPP 052 v1.1 (July 7, 1996)
    -- Taps are 1-based such that zero denotes the tap is not required.
    constant C_TAPTABLE : t_taptable := (
        (  3,   2,   0,   0,   0), --   3
        (  4,   3,   0,   0,   0), --   4
        (  5,   3,   0,   0,   0), --   5
        (  6,   5,   0,   0,   0), --   6
        (  7,   6,   0,   0,   0), --   7
        (  8,   6,   5,   4,   0), --   8
        (  9,   5,   0,   0,   0), --   9
        ( 10,   7,   0,   0,   0), --  10
        ( 11,   9,   0,   0,   0), --  11
        ( 12,   6,   4,   1,   0), --  12
        ( 13,   4,   3,   1,   0), --  13
        ( 14,   5,   3,   1,   0), --  14
        ( 15,  14,   0,   0,   0), --  15
        ( 16,  15,  13,   4,   0), --  16
        ( 17,  14,   0,   0,   0), --  17
        ( 18,  11,   0,   0,   0), --  18
        ( 19,   6,   2,   1,   0), --  19
        ( 20,  17,   0,   0,   0), --  20
        ( 21,  19,   0,   0,   0), --  21
        ( 22,  21,   0,   0,   0), --  22
        ( 23,  18,   0,   0,   0), --  23
        ( 24,  23,  22,  17,   0), --  24
        ( 25,  22,   0,   0,   0), --  25
        ( 26,   6,   2,   1,   0), --  26
        ( 27,   5,   2,   1,   0), --  27
        ( 28,  25,   0,   0,   0), --  28
        ( 29,  27,   0,   0,   0), --  29
        ( 30,   6,   4,   1,   0), --  30
        ( 31,  28,   0,   0,   0), --  31
        ( 32,  22,   2,   1,   0), --  32
        ( 33,  20,   0,   0,   0), --  33
        ( 34,  27,   2,   1,   0), --  34
        ( 35,  33,   0,   0,   0), --  35
        ( 36,  25,   0,   0,   0), --  36
        ( 37,   5,   4,   3,   2), --  37
        ( 38,   6,   5,   1,   0), --  38
        ( 39,  35,   0,   0,   0), --  39
        ( 40,  38,  21,  19,   0), --  40
        ( 41,  38,   0,   0,   0), --  41
        ( 42,  41,  20,  19,   0), --  42
        ( 43,  42,  38,  37,   0), --  43
        ( 44,  43,  18,  17,   0), --  44
        ( 45,  44,  42,  41,   0), --  45
        ( 46,  45,  26,  25,   0), --  46
        ( 47,  42,   0,   0,   0), --  47
        ( 48,  47,  21,  20,   0), --  48
        ( 49,  40,   0,   0,   0), --  49
        ( 50,  49,  24,  23,   0), --  50
        ( 51,  50,  36,  35,   0), --  51
        ( 52,  49,   0,   0,   0), --  52
        ( 53,  52,  38,  37,   0), --  53
        ( 54,  53,  18,  17,   0), --  54
        ( 55,  31,   0,   0,   0), --  55
        ( 56,  55,  35,  34,   0), --  56
        ( 57,  50,   0,   0,   0), --  57
        ( 58,  39,   0,   0,   0), --  58
        ( 59,  58,  38,  37,   0), --  59
        ( 60,  59,   0,   0,   0), --  60
        ( 61,  60,  46,  45,   0), --  61
        ( 62,  61,   6,   5,   0), --  62
        ( 63,  62,   0,   0,   0), --  63
        ( 64,  63,  61,  60,   0), --  64
        ( 65,  47,   0,   0,   0), --  65
        ( 66,  65,  57,  56,   0), --  66
        ( 67,  66,  58,  57,   0), --  67
        ( 68,  59,   0,   0,   0), --  68
        ( 69,  67,  42,  40,   0), --  69
        ( 70,  69,  55,  54,   0), --  70
        ( 71,  65,   0,   0,   0), --  71
        ( 72,  66,  25,  19,   0), --  72
        ( 73,  48,   0,   0,   0), --  73
        ( 74,  73,  59,  58,   0), --  74
        ( 75,  74,  65,  64,   0), --  75
        ( 76,  75,  41,  40,   0), --  76
        ( 77,  76,  47,  46,   0), --  77
        ( 78,  77,  59,  58,   0), --  78
        ( 79,  70,   0,   0,   0), --  79
        ( 80,  79,  43,  42,   0), --  80
        ( 81,  77,   0,   0,   0), --  81
        ( 82,  79,  47,  44,   0), --  82
        ( 83,  82,  38,  37,   0), --  83
        ( 84,  71,   0,   0,   0), --  84
        ( 85,  84,  58,  57,   0), --  85
        ( 86,  85,  74,  73,   0), --  86
        ( 87,  74,   0,   0,   0), --  87
        ( 88,  87,  17,  16,   0), --  88
        ( 89,  51,   0,   0,   0), --  89
        ( 90,  89,  72,  71,   0), --  90
        ( 91,  90,   8,   7,   0), --  91
        ( 92,  91,  80,  79,   0), --  92
        ( 93,  91,   0,   0,   0), --  93
        ( 94,  73,   0,   0,   0), --  94
        ( 95,  84,   0,   0,   0), --  95
        ( 96,  94,  49,  47,   0), --  96
        ( 97,  91,   0,   0,   0), --  97
        ( 98,  87,   0,   0,   0), --  98
        ( 99,  97,  54,  52,   0), --  99
        (100,  63,   0,   0,   0), -- 100
        (101, 100,  95,  94,   0), -- 101
        (102, 101,  36,  35,   0), -- 102
        (103,  94,   0,   0,   0), -- 103
        (104, 103,  94,  93,   0), -- 104
        (105,  89,   0,   0,   0), -- 105
        (106,  91,   0,   0,   0), -- 106
        (107, 105,  44,  42,   0), -- 107
        (108,  77,   0,   0,   0), -- 108
        (109, 108, 103, 102,   0), -- 109
        (110, 109,  98,  97,   0), -- 110
        (111, 101,   0,   0,   0), -- 111
        (112, 110,  69,  67,   0), -- 112
        (113, 104,   0,   0,   0), -- 113
        (114, 113,  33,  32,   0), -- 114
        (115, 114, 101, 100,   0), -- 115
        (116, 115,  46,  45,   0), -- 116
        (117, 115,  99,  97,   0), -- 117
        (118,  85,   0,   0,   0), -- 118
        (119, 111,   0,   0,   0), -- 119
        (120, 113,   9,   2,   0), -- 120
        (121, 103,   0,   0,   0), -- 121
        (122, 121,  63,  62,   0), -- 122
        (123, 121,   0,   0,   0), -- 123
        (124,  87,   0,   0,   0), -- 124
        (125, 124,  18,  17,   0), -- 125
        (126, 125,  90,  89,   0), -- 126
        (127, 126,   0,   0,   0), -- 127
        (128, 126, 101,  99,   0), -- 128
        (129, 124,   0,   0,   0), -- 129
        (130, 127,   0,   0,   0), -- 130
        (131, 130,  84,  83,   0), -- 131
        (132, 103,   0,   0,   0), -- 132
        (133, 132,  82,  81,   0), -- 133
        (134,  77,   0,   0,   0), -- 134
        (135, 124,   0,   0,   0), -- 135
        (136, 135,  11,  10,   0), -- 136
        (137, 116,   0,   0,   0), -- 137
        (138, 137, 131, 130,   0), -- 138
        (139, 136, 134, 131,   0), -- 139
        (140, 111,   0,   0,   0), -- 140
        (141, 140, 110, 109,   0), -- 141
        (142, 121,   0,   0,   0), -- 142
        (143, 142, 123, 122,   0), -- 143
        (144, 143,  75,  74,   0), -- 144
        (145,  93,   0,   0,   0), -- 145
        (146, 145,  87,  86,   0), -- 146
        (147, 146, 110, 109,   0), -- 147
        (148, 121,   0,   0,   0), -- 148
        (149, 148,  40,  39,   0), -- 149
        (150,  97,   0,   0,   0), -- 150
        (151, 148,   0,   0,   0), -- 151
        (152, 151,  87,  86,   0), -- 152
        (153, 152,   0,   0,   0), -- 153
        (154, 152,  27,  25,   0), -- 154
        (155, 154, 124, 123,   0), -- 155
        (156, 155,  41,  40,   0), -- 156
        (157, 156, 131, 130,   0), -- 157
        (158, 157, 132, 131,   0), -- 158
        (159, 128,   0,   0,   0), -- 159
        (160, 159, 142, 141,   0), -- 160
        (161, 143,   0,   0,   0), -- 161
        (162, 161,  75,  74,   0), -- 162
        (163, 162, 104, 103,   0), -- 163
        (164, 163, 151, 150,   0), -- 164
        (165, 164, 135, 134,   0), -- 165
        (166, 165, 128, 127,   0), -- 166
        (167, 161,   0,   0,   0), -- 167
        (168, 166, 153, 151,   0)  -- 168
    );

    ----------------------------------------------------------------------------
    -- Procedure: LFSR Advance
    -- * Advances LFSR register by one.
    -- * Size is inferred from the input arguments.
    ----------------------------------------------------------------------------
    procedure lfsr_advance (
        signal REG : inout std_logic_vector
    );

    ----------------------------------------------------------------------------
    -- Procedure: LFSR Advance
    -- * Advances LFSR register by one, up to a desired reset value.
    -- * LFSR resets after the reset value is reached.
    -- * Size is inferred from the input arguments.
    ----------------------------------------------------------------------------
    procedure lfsr_advance (
        signal REG : inout std_logic_vector;
        constant RESET : in std_logic_vector
    );

    ----------------------------------------------------------------------------
    -- Procedure: LFSR Advance (Variable)
    -- * Advances LFSR variable by one.
    -- * Size is inferred from the input arguments.
    ----------------------------------------------------------------------------
    procedure lfsr_advance_var (
        variable REG : inout std_logic_vector
    );

    ----------------------------------------------------------------------------
    -- Procedure: LFSR Advance (Variable)
    -- * Advances LFSR variable by one, up to a desired reset value.
    -- * LFSR resets after the reset value is reached.
    -- * Size is inferred from the input arguments.
    ----------------------------------------------------------------------------
    procedure lfsr_advance_var (
        variable REG : inout std_logic_vector;
        constant RESET : in std_logic_vector
    );

    ----------------------------------------------------------------------------
    -- Function: LFSR Evaluate
    -- * Calculate the LFSR register value reached after a chosen number of
    --   iterations.
    -- * Size must be given as it cannot be inferred from the input arguments.
    ----------------------------------------------------------------------------
    function lfsr_evaluate (
        constant SIZE : natural;
        constant VALUE : natural
    ) return std_logic_vector;

    ----------------------------------------------------------------------------
    -- Function: LFSR Maximum
    -- * Calculate the maximum sequence length for a chosen LFSR size.
    -- * Size must be given as it cannot be inferred from the input arguments.
    ----------------------------------------------------------------------------
    function lfsr_maximum (constant SIZE : natural) return natural;

end lfsr;
--------------------------------------------------------------------------------